magic
tech sky130A
timestamp 1720323565
<< nwell >>
rect -350 0 -50 380
<< nmos >>
rect -210 -250 -195 -100
<< pmos >>
rect -210 50 -195 250
<< ndiff >>
rect -300 -115 -210 -100
rect -300 -235 -285 -115
rect -230 -235 -210 -115
rect -300 -250 -210 -235
rect -195 -115 -105 -100
rect -195 -235 -175 -115
rect -120 -235 -105 -115
rect -195 -250 -105 -235
<< pdiff >>
rect -300 235 -210 250
rect -300 65 -285 235
rect -230 65 -210 235
rect -300 50 -210 65
rect -195 235 -105 250
rect -195 65 -175 235
rect -120 65 -105 235
rect -195 50 -105 65
<< ndiffc >>
rect -285 -235 -230 -115
rect -175 -235 -120 -115
<< pdiffc >>
rect -285 65 -230 235
rect -175 65 -120 235
<< psubdiff >>
rect -300 -310 -100 -290
rect -300 -330 -270 -310
rect -130 -330 -100 -310
rect -300 -345 -100 -330
<< nsubdiff >>
rect -300 335 -100 350
rect -300 315 -275 335
rect -125 315 -100 335
rect -300 300 -100 315
<< psubdiffcont >>
rect -270 -330 -130 -310
<< nsubdiffcont >>
rect -275 315 -125 335
<< poly >>
rect -210 250 -195 265
rect -210 -10 -195 50
rect -285 -25 -195 -10
rect -285 -50 -265 -25
rect -240 -50 -195 -25
rect -285 -65 -195 -50
rect -210 -100 -195 -65
rect -210 -265 -195 -250
<< polycont >>
rect -265 -50 -240 -25
<< locali >>
rect -300 335 -100 350
rect -300 315 -275 335
rect -125 315 -100 335
rect -300 300 -100 315
rect -300 250 -235 300
rect -300 235 -215 250
rect -300 65 -285 235
rect -230 65 -215 235
rect -300 50 -215 65
rect -190 235 -105 250
rect -190 65 -175 235
rect -120 65 -105 235
rect -190 50 -105 65
rect -345 -25 -215 -10
rect -345 -50 -310 -25
rect -290 -50 -265 -25
rect -240 -50 -215 -25
rect -345 -65 -215 -50
rect -170 -30 -105 50
rect -170 -55 -145 -30
rect -125 -55 -105 -30
rect -170 -100 -105 -55
rect -300 -115 -215 -100
rect -300 -235 -285 -115
rect -230 -235 -215 -115
rect -300 -250 -215 -235
rect -190 -115 -105 -100
rect -190 -235 -175 -115
rect -120 -235 -105 -115
rect -190 -250 -105 -235
rect -295 -295 -230 -250
rect -295 -310 -105 -295
rect -295 -330 -270 -310
rect -130 -330 -105 -310
rect -295 -340 -105 -330
<< viali >>
rect -245 315 -160 335
rect -310 -50 -290 -25
rect -145 -55 -125 -30
rect -245 -330 -145 -310
<< metal1 >>
rect -345 335 -55 350
rect -345 315 -245 335
rect -160 315 -55 335
rect -345 300 -55 315
rect -350 -25 -270 -10
rect -350 -50 -310 -25
rect -290 -50 -270 -25
rect -350 -65 -270 -50
rect -160 -30 20 -10
rect -160 -55 -145 -30
rect -125 -55 20 -30
rect -160 -70 20 -55
rect -350 -310 -55 -290
rect -350 -330 -245 -310
rect -145 -330 -55 -310
rect -350 -345 -55 -330
<< labels >>
rlabel metal1 -350 -55 -350 -55 3 vin
rlabel metal1 -45 -50 -45 -50 1 vout
rlabel metal1 -75 -330 -75 -330 1 vss
rlabel metal1 -80 325 -80 325 1 vdd
<< end >>
